Vim�UnDo� /�f��J1�-�)��Q�(�M���`�6�   `   module uart(            �       �   �   �    `>)�   � _�                             ����                                                                                                                                                                                                                                                                                                                                                             `<�    �                R//////////////////////////////////////////////////////////////////////////////////   // Company:    // Engineer:    //    #// Create Date: 2021/03/01 21:40:48   // Design Name:    // Module Name: uart   // Project Name:    // Target Devices:    // Tool Versions:    // Description:    //    // Dependencies:    //    // Revision:   // Revision 0.01 - File Created   // Additional Comments:   //    R//////////////////////////////////////////////////////////////////////////////////5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `<�%    �                5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `<��     �         	      		input sys_clk,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `<��    �         	      		input sys_rst_n,5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `=�    �                		5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `=�    �      	         	input sys_rst_n,   );�                   );5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `=�     �      	   	    5�_�      	                      ����                                                                                                                                                                                                                                                                                                                                                             `=�    �      
   	       5�_�      
           	   	       ����                                                                                                                                                                                                                                                                                                                                                             `=�Q     �   	   
       5�_�   	              
   	       ����                                                                                                                                                                                                                                                                                                                                                             `=�Z    �      
         	output uart_date,5�_�   
                 	       ����                                                                                                                                                                                                                                                                                                                                                             `=�d     �   	   
       5�_�                    	       ����                                                                                                                                                                                                                                                                                                                                                             `=�f    �   	            	�   	          5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             `=�w   
 �   
          5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `=��    �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `=��    �             5�_�                    
       ����                                                                                                                                                                                                                                                                                                                                                             `=��    �   	            	output uart_done,5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `>X    �                5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `>`     �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `>b    �                5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               	reg urat_rxd0,uart_rxd1;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               	reg urat_rxd0uart_rxd1;5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               	reg urat_rxd05�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�                       
    ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               		uart_rxd15�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               		uart_rxd05�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             `>�    �             5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             `>�    �             5�_�      !                     ����                                                                                                                                                                                                                                                                                                                                                             `>�    �               		�             5�_�      "           !           ����                                                                                                                                                                                                                                                                                                                                                             `>-    �                 5�_�   !   #           "      	    ����                                                                                                                                                                                                                                                                                                                                                             `>4    �               			if(!sys5�_�   "   $           #          ����                                                                                                                                                                                                                                                                                                                                                             `>H    �             5�_�   #   %           $          ����                                                                                                                                                                                                                                                                                                                                                             `>N    �               		uart_rxd0<=1'b1;5�_�   $   &           %          ����                                                                                                                                                                                                                                                                                                                                                             `>O     �             5�_�   %   '           &           ����                                                                                                                                                                                                                                                                                                                                                             `>T     �                5�_�   &   (           '          ����                                                                                                                                                                                                                                                                                                                                                             `>W     �             5�_�   '   )           (          ����                                                                                                                                                                                                                                                                                                                                                             `>Y   ! �               		�             5�_�   (   *           )          ����                                                                                                                                                                                                                                                                                                                                                             `>]   " �             5�_�   )   +           *          ����                                                                                                                                                                                                                                                                                                                                                             `>k   # �               	reg urat_rxd0;5�_�   *   ,           +          ����                                                                                                                                                                                                                                                                                                                                                             `>l   $ �               	reg urt_rxd0;5�_�   +   -           ,          ����                                                                                                                                                                                                                                                                                                                                                             `>n   % �               	reg ur_rxd0;5�_�   ,   .           -          ����                                                                                                                                                                                                                                                                                                                                                             `>s   & �               	reg u_rxd0;5�_�   -   1           .          ����                                                                                                                                                                                                                                                                                                                                                             `>u   ) �             5�_�   .   2   /       1          ����                                                                                                                                                                                                                                                                                                                                                             `>�   * �               			�             5�_�   1   3           2          ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                                                             `>�   + �               		�             5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                                                             `>�   , �             5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                                                             `>   - �               	�             5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                                                             `>     �             5�_�   6   8           7          ����                                                                                                                                                                                                                                                                                                                                                             `>   . �               	�             5�_�   7   9           8          ����                                                                                                                                                                                                                                                                                                                                                             `>.     �             5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                             `>�   / �               	assign 5�_�   9   ;           :      (    ����                                                                                                                                                                                                                                                                                                                                                             `>�   0 �             5�_�   :   <           ;          ����                                                                                                                                                                                                                                                                                                                                                             `>   1 �               *	assign start_flag=uart_rxd1(~uart_rxd0); 5�_�   ;   =           <          ����                                                                                                                                                                                                                                                                                                                                                             `>   2 �             5�_�   <   >           =          ����                                                                                                                                                                                                                                                                                                                                                             `>{   3 �               	�             5�_�   =   ?           >          ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�   >   @           ?          ����                                                                                                                                                                                                                                                                                                                                                             `>�   4 �               	reg 5�_�   ?   A           @          ����                                                                                                                                                                                                                                                                                                                                                             `>�   5 �             5�_�   @   B           A           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   6 �                �             5�_�   A   C           B      2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   7 �      $         2	always @(posedge sys_clk,negedge sys_rst_n) begin5�_�   B   D           C   #       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�     �   #   $   $    5�_�   C   E           D          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   8 �         $      		if(!sys_rst_n) begin5�_�   D   F           E          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>     �         $    5�_�   E   G           F            ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   9 �      !   $       5�_�   F   H           G           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>'     �       !   $    5�_�   G   I           H           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>+   : �                 5�_�   H   J           I           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>,   ; �                 		end5�_�   I   K           J          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>1   < �         "      		if(!sys_rst_n) begin5�_�   J   L           K          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>2   = �         "      		if(!sys_rst_n) egin5�_�   K   M           L          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>2   > �         "      		if(!sys_rst_n) gin5�_�   L   N           M          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>2   ? �         "      		if(!sys_rst_n) in5�_�   M   O           N          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>2   @ �         "      		if(!sys_rst_n) n5�_�   N   P           O            ����                                                                                                                                                                                                                                                                                                                               1                  v        `>8   A �      !   "       5�_�   O   S           P           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>a   C �       !   "    5�_�   P   T   Q       S          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>k   D �         #      	�         "    5�_�   S   U           T           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>     �         %    5�_�   T   V           U   #       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   E �   "   &   %      		else 5�_�   U   W           V   %   #    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�     �   %   &   '    5�_�   V   X           W           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   F �         (      	�         '    5�_�   W   Y           X           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   G �         +    5�_�   X   Z           Y   )   $    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   H �   (   *   +      $		else if(rx_cnt==4'd9)&&(clk_cnt ==5�_�   Y   [           Z   )   1    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   I �   )   *   +    5�_�   Z   \           [   )   1    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>-   J �   )   ,   ,      			�   )   +   +    5�_�   [   ]           \   +       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>J     �   +   ,   -    5�_�   \   ^           ]   *       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>K   K �   )   +   -      			rx_flag<=1'b1;5�_�   ]   _           ^   *       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>O   L �   )   +   -      			rx_flag<=1'b;5�_�   ^   `           _   *       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>P     �   *   +   -    5�_�   _   a           `   +       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>T   M �   *   ,   -      		5�_�   `   b           a   +       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>     �   +   ,   -    5�_�   a   c           b   +       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   N �   *   ,   -      			u5�_�   b   d           c   )   2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   O �   (   *   -      2		else if(rx_cnt==4'd9)&&(clk_cnt == BPS_CNT-1'b1)5�_�   c   e           d   )   2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   P �   )   *   -    5�_�   d   f           e   )   2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   Q �   (   *   -      3		else if(rx_cnt==4'd9)&&(clk_cnt == BPS_CNT-1'b1);5�_�   e   g           f   )   2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   R �   (   *   -      2		else if(rx_cnt==4'd9)&&(clk_cnt == BPS_CNT-1'b1)5�_�   f   h           g   )   2    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�     �   )   *   -    5�_�   g   i           h   )   	    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�   S �   (   *   -      3		else if(rx_cnt==4'd9)&&(clk_cnt == BPS_CNT-1'b1))5�_�   h   j           i   )   	    ����                                                                                                                                                                                                                                                                                                                               1                  v        `>�     �   )   *   -    5�_�   i   k           j   ,       ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   T �   ,   .   -    5�_�   j   n           k   -        ����                                                                                                                                                                                                                                                                                                                               1                  v        `>   X �   -   .   .    5�_�   k   o   m       n   -        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>$   Y �   ,   0   .       �   -   .   .    5�_�   n   p           o   /        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>)   Z �   /   1   1      			�   /   1   0    5�_�   o   q           p   0       ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>-     �   0   1   1    5�_�   p   r           q   /        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>7   [ �   -   2   1      		if(!sys_rst_n)     �   .   0   1       5�_�   q   s           r   1        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>z     �   1   2   3    5�_�   r   t           s   1        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>�   \ �   /   4   3      		else if(rx_flag) begin    �   0   2   3       5�_�   s   u           t   3       ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>�     �   3   4   5    5�_�   t   v           u   0       ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>�   ] �   0   6   6      			�   0   2   5    5�_�   u   w           v   5        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>�   ^ �   5   6   :    5�_�   v   x           w   5        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	   _ �   4   5           5�_�   w   y           x   8       ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	   ` �   8   :   9    5�_�   x   z           y   9        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>		     �   9   :   :    5�_�   y   {           z   9        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	
   a �   9   ;   :    �   9   :   :    5�_�   z   |           {   9        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	   b �   8   <   ;       �   9   :   ;    5�_�   {   }           |   ;        ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	&   c �   :   @   =       5�_�   |   ~           }   ?       ����                                                                                                                                                                                                                                                                                                                            $           %          v���    `>	?   e �   ?   @   A    5�_�   }              ~   =        ����                                                                                                                                                                                                                                                                                                                            #           A           v        `> �   f �   <   =           5�_�   ~   �              <       ����                                                                                                                                                                                                                                                                                                                            #           @           v        `> �   g �   ;   B   @      		else5�_�      �           �   A       ����                                                                                                                                                                                                                                                                                                                            #           E           v        `>!     �   A   B   E    5�_�   �   �           �   B        ����                                                                                                                                                                                                                                                                                                                            #           E           v        `>!   h �   A   B           5�_�   �   �           �   A       ����                                                                                                                                                                                                                                                                                                                            #           D           v        `>!   i �   @   B   D      			5�_�   �   �           �   A       ����                                                                                                                                                                                                                                                                                                                            #           D           v        `>!     �   A   B   D    5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                            #           D           v        `>!'   j �         D       5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                            #           D           v        `>!3     �         D    5�_�   �   �           �   C        ����                                                                                                                                                                                                                                                                                                                            #           D           v        `>!:   k �   C   E   D    �   C   D   D    5�_�   �   �           �   C        ����                                                                                                                                                                                                                                                                                                                            #           E           v        `>!>   l �   B   F   E       �   C   D   E    5�_�   �   �           �   E        ����                                                                                                                                                                                                                                                                                                                            #           G           v        `>!E     �   C   J   G      		if(!sys_rst_n)     �   D   F   G       5�_�   �   �           �   H        ����                                                                                                                                                                                                                                                                                                                            #           K           v        `>!�   m �   G   J   K       5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                            #           L           v        `>"+     �   I   J   L    5�_�   �   �           �   F       ����                                                                                                                                                                                                                                                                                                                            #           L           v        `>"8   n �   E   G   L      		else if(rx_flag) begin5�_�   �   �           �   F   &    ����                                                                                                                                                                                                                                                                                                                            #           L           v        `>"W   q �   F   G   L    5�_�   �   �   �       �   I        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"r   r �   H   K   L       �   I   J   L    5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"r   s �   H   K   M      				4'd1:rxdata[0]<=uart_rxd1;�   I   J   M    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"s   t �   H   K   N      					4'd1:rxdata[0]<=uart_rxd1;�   I   J   N    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"s   u �   H   K   O       						4'd1:rxdata[0]<=uart_rxd1;�   I   J   O    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"t   v �   H   K   P      !							4'd1:rxdata[0]<=uart_rxd1;�   I   J   P    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"u   w �   H   K   Q      "								4'd1:rxdata[0]<=uart_rxd1;�   I   J   Q    5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"x   x �   H   J   R      #									4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"x   y �   H   J   R      "								4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"x   z �   H   J   R      !							4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"y   { �   H   J   R       						4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"|   | �   H   J   R      					4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"|   } �   H   J   R      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   H   J   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   I   K   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   J   L   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   K   M   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   L   N   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   ~ �   M   O   R      			4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�     �   N   O   R    5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�    �   N   P   R       �   O   P   R    5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   N   Q   R      	�   O   P   R    5�_�   �   �           �   O        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   N   P   S      					4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   H   J   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   I   K   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   J   L   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   K   M   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   L   N   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   M   O   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   N   P   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   H   J   S      				4'd2:rxdata[0]<=uart_rxd1;5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   I   K   S      				4'd3:rxdata[0]<=uart_rxd1;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   J   L   S      				4'd4:rxdata[0]<=uart_rxd1;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   K   M   S      				4'd5:rxdata[0]<=uart_rxd1;5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   L   N   S      				4'd6:rxdata[0]<=uart_rxd1;5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   M   O   S      				4'd7:rxdata[0]<=uart_rxd1;5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   N   P   S      				4'd8:rxdata[0]<=uart_rxd1;5�_�   �   �   �       �   R        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   Q   S   S       5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   R   S   S    5�_�   �   �           �   R       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   R   T   T      		�   R   T   S    5�_�   �   �           �   S       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   S   T   T    5�_�   �   �           �   P        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   O   P           5�_�   �   �           �   H       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   G   I   S      				4'd1:rxdata[0]<=uart_rxd1;5�_�   �   �           �   I       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   H   J   S      				4'd2:rxdata[1]<=uart_rxd1;5�_�   �   �           �   J       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   I   K   S      				4'd3:rxdata[2]<=uart_rxd1;5�_�   �   �           �   K       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   J   L   S      				4'd4:rxdata[3]<=uart_rxd1;5�_�   �   �           �   L       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   K   M   S      				4'd5:rxdata[4]<=uart_rxd1;5�_�   �   �           �   M       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   L   N   S      				4'd6:rxdata[5]<=uart_rxd1;5�_�   �   �           �   N       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#     �   M   O   S      				4'd7:rxdata[6]<=uart_rxd1;5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#   � �   N   P   S      				4'd8:rxdata[7]<=uart_rxd1;5�_�   �   �           �   O       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#   � �   O   P   S    5�_�   �   �           �   R        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#\   � �   R   T   S    5�_�   �   �           �   S        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#\     �   S   T   T    5�_�   �   �           �   S        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#b   � �   R   V   T       �   S   T   T    5�_�   �   �           �   T        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#f     �   T   V   W      			�   T   V   V    5�_�   �   �           �   V        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#n     �   U   W   W       5�_�   �   �           �   U       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#u   � �   S   Z   W      		if(!sys_rst_n)    	�   T   V   W      		5�_�   �   �           �   Y        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�     �   Y   Z   [    5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�   � �      
   [      	output [7:0] uart_date,5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�     �   	   
   [    5�_�   �   �           �   
       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�   � �   	      [      	output uart_done5�_�   �   �           �   
       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�     �   
      [    5�_�   �   �           �   X       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>#�   � �   W   _   [      		else5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$L     �   ^   _   a    5�_�   �   �           �   \        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$�   � �   [   \           5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$�   � �   \   _   `      			uart_data5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$�     �   ^   _   a    5�_�   �   �           �   ]       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$�   � �   \   ^   a      			uart_data<=1'b0;5�_�   �   �           �   _        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>$�   � �   ^   `   a       5�_�   �   �           �   _       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%      �   _   `   a    5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%   � �   ]   _   a      			urat_done<=1'b0;5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%   � �   ]   _   a      			uat_done<=1'b0;5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%   � �   ]   _   a      			ut_done<=1'b0;5�_�   �   �           �   ^       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%     �   ^   _   a    5�_�   �   �           �   	       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%P   � �      
   a      	output reg [7:0] uart_date,5�_�   �   �           �   V       ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>%[   � �   U   W   a      			uart_date<=8'b0;5�_�   �   �           �   )   -    ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>&   � �   (   *   a      4		else if((rx_cnt==4'd9)&&(clk_cnt == BPS_CNT-1'b1))5�_�   �   �   �       �           ����                                                                                                                                                                                                                                                                                                                                                             `>)z   � �                    module uart(   	input sys_clk,   	input sys_rst_n,   	   	input uart_rxd,   	output [7:0] uart_date,   	output uart_done   );   	reg urat_rxd0;   	reg uart_rxd1;   2	always @(posedge sys_clk,negedge sys_rst_n) begin   		uart_rxd0<=1'b1;           	endmodule5�_�   �   �           �           ����                                                                                                                                                                                                                                                                                                                                                             `>)   � �                  �               5�_�   �   �           �          ����                                                                                                                                                                                                                                                                                                                                                             `>)�   � �         `      module uart(5�_�   �               �          ����                                                                                                                                                                                                                                                                                                                                                             `>)�   � �         `    5�_�   �           �   �   )   .    ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>&   � �   )   *   a    5�_�   �           �   �   R        ����                                                                                                                                                                                                                                                                                                                            H           H          v���    `>"�   � �   Q   T        5�_�   �           �   �   I        ����                                                                                                                                                                                                                                                                                                                            H          H          v���    `>"i   p �   I   J   L    �   H   J   L      4'd1:rxdata[0]<=uart_rxd1;    5�_�   k       l   n   m   $        ����                                                                                                                                                                                                                                                                                                                            $           $           v���    `>   W �   #   '   .      		rx_flag<=1'b0;�   $   %   ,    �   #   %   ,      ;		rx_flag<=1'b0;5�_�   k           m   l   -        ����                                                                                                                                                                                                                                                                                                                               1                  v        `>
   U �   -   .   .    �   ,   .   .      ;;;;5�_�   P   R       S   Q          ����                                                                                                                                                                                                                                                                                                                               1                  v        `>g   B �         "       5�_�   Q               R           ����                                                                                                                                                                                                                                                                                                                               1                  v        `>h     �         #    5�_�   .   0       1   /          ����                                                                                                                                                                                                                                                                                                                                                             `>�   ( �                5�_�   /               0           ����                                                                                                                                                                                                                                                                                                                                                             `>�     �             5�_�              !               ����                                                                                                                                                                                                                                                                                                                                                             `>     �             5��